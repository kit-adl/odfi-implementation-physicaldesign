VERSION 5.6 ;

MACRO ExampleMacro_333x105
  CLASS BLOCK ; 
  ORIGIN 0 0 ;
  SIZE 333.42 BY 105.28 ;
END ExampleMacro_333x105

MACRO ExampleMacro_50x50
  CLASS BLOCK ; 
  ORIGIN 0 0 ;
  SIZE 50 BY 50 ;
END ExampleMacro_50x50

END LIBRARY
